library verilog;
use verilog.vl_types.all;
entity counter6_vlg_sample_tst is
    port(
        cp              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end counter6_vlg_sample_tst;
