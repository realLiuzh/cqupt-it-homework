library verilog;
use verilog.vl_types.all;
entity code_select_vlg_check_tst is
    port(
        t_04            : in     vl_logic_vector(3 downto 0);
        sampler_rx      : in     vl_logic
    );
end code_select_vlg_check_tst;
