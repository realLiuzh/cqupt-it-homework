library verilog;
use verilog.vl_types.all;
entity counter6_vlg_vec_tst is
end counter6_vlg_vec_tst;
